`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/11/18 16:27:11
// Design Name: 
// Module Name: half_adder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module half_adder(
input a,input b, 
output sum,output c_out
); //�����
     //xor �޽�λ�ӷ�
     assign sum = a^b;
     //��λ��Ϣ1&1=1����λ
     assign c_out = a&b;
endmodule
